* AC Analysis, 500 lowPass, 9th order Chebyshev 3 dB, 5 stages using AD8617

* Input signal for AC and transient sinusoidal analysis 
VIN IN 0 AC 1 DC 2.5 SIN(2.5 1.59 50) 
* VNOISE IN 0 AC 0 DC 2.5 

XA IN OUTA VCCG VEEG 0 firstOrderlowPassStageA
XB OUTA OUTB VCCG VEEG 0 sallenKeylowPassStageB
XC OUTB OUTC VCCG VEEG 0 sallenKeylowPassStageC
XD OUTC OUTD VCCG VEEG 0 sallenKeylowPassStageD
XE OUTD OUT VCCG VEEG 0 sallenKeylowPassStageE

VP VCCG 0 5
VM VEEG 0 0

*Simulation directive lines for AC Analysis 
.AC DEC 100 50 6E3 
*.TRAN 1ns 7.98E-3 
*.NOISE V(OUT) VNOISE DEC 100 50 6E3 
.PROBE 

.SUBCKT firstOrderlowPassStageA IN OUT VCC VEE GND 
X1 INP OUT VCC VEE OUT AD8617 
R1 IN INP 98.2E3 
C1 INP GND 33E-9 
.ENDS firstOrderlowPassStageA 

.SUBCKT sallenKeylowPassStageB IN OUT VCC VEE GND 
X1 INP OUT VCC VEE OUT AD8617 
R1 IN 1 379E3 
R2 1 INP 379E3 
C1 1 OUT 9.1E-9 
C2 INP GND 613E-12 
.ENDS sallenKeylowPassStageB 

.SUBCKT sallenKeylowPassStageC IN OUT VCC VEE GND 
X1 INP OUT VCC VEE OUT AD8617 
R1 IN 1 46.5E3 
R2 1 INP 46.5E3 
C1 1 OUT 91E-9 
C2 INP GND 1.22E-9 
.ENDS sallenKeylowPassStageC 

.SUBCKT sallenKeylowPassStageD IN OUT VCC VEE GND 
X1 INP OUT VCC VEE OUT AD8617 
R1 IN 1 5.4E3 
R2 1 INP 5.4E3 
C1 1 OUT 1.2E-6 
C2 INP GND 3.81E-9 
.ENDS sallenKeylowPassStageD 

.SUBCKT sallenKeylowPassStageE IN OUT VCC VEE GND 
X1 INP OUT VCC VEE OUT AD8617 
R1 IN 1 20.5E3 
R2 1 INP 20.5E3 
C1 1 OUT 910E-9 
C2 INP GND 271E-12 
.ENDS sallenKeylowPassStageE 

* AD8617 SPICE Macro-model
* Description: Amplifier
* Generic Desc: 1.8/5V, CMOS, OP, Low Pwr, RRIO, 2X
* Developed by: VW ADSJ
* Revision History: 08/10/2012 - Updated to new header style
* 2.0 (02/2010)
* 3.0 (03/2017) - Followed AD8613 model, dual version only
* Copyright 2010, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes: VSY=5V, T=25degC
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8617          1   2   99  50  45
*#ASSOC Category="Op-amps" symbol=opamp
*
* INPUT STAGE
*
M1  14  7  8  8 PIX L=1E-6 W=2.37E-04
M2  16  2  8  8 PIX L=1E-6 W=2.37E-04
M3  17  7 10 10 NIX L=1E-6 W=8.88E-05
M4  18  2 10 10 NIX L=1E-6 W=8.88E-05
RD1 14 50 8.00E+04
RD2 16 50 8.00E+04
RD3 99 17 8.00E+04
RD4 99 18 8.00E+04
C1  14 16 8.08E-13
C2  17 18 8.08E-13
I1  99  8 5.00E-06
I2  10 50 5.00E-06
V1  99  9 2.625E-01
V2  13 50 1.625E-01
D1   8  9 DX
D2  13 10 DX
EOS  7  1 POLY(4) (22,98) (73,98) (81,98) (70,98) 4.00E-04 1 1 1 1
IOS  1  2 5.00E-14
*
*CMRR=95dB, POLE AT 1000 Hz
*
E1  21 98 POLY(2) (1,98) (2,98) 0 8.89E-03 8.89E-03
R10 21 22 1.59E+04
R20 22 98 1.59E-01
C10 21 22 1.00E-09
*
* PSRR=90dB, POLE AT 100 Hz
*
EPSY 72 98 POLY(1) (99,50) -1.58113883 0.316227766
CPS3 72 73 1.00E-06
RPS3 72 73 1.59E+03
RPS4 73 98 1.59E-01
*
* VOLTAGE NOISE REFERENCE OF 22nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 1.98E+01
RN2 81 98 1
*
* FLICKER NOISE CORNER = 100 Hz
*
D5  69 98 DNOISE
VSN 69 98 DC 0.6551
H1  70 98 POLY(1) VSN 1.00E-03 1.00E+00
RN  70 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) -8.09E-06 3.0E-06
EVP  97 98 POLY(1) (99,50) 0 0.5
EVN  51 98 POLY(1) (50,99) 0 0.5
*
* GAIN STAGE
*
G1 98 30 POLY(2) (14,16) (17,18) 0 4.15E-05 4.15E-05
R1 30 98 1.00E+06
RZ 30 31 7.91E+02
CF 45 31 3.32E-10
V3 32 30 3.53E-01
V4 30 33 -7.53E-01
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=1E-6 W=2.50E-04
M6  45 47 50 50 NOX L=1E-6 W=1.93E-03
EG1 99 46 POLY(1) (98,30) 7.465E-01 1
EG2 47 50 POLY(1) (30,98) 6.335E-01 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=4.00E-05,VTO=-0.7,LAMBDA=0.047,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=1.00E-05,VTO=+0.6,LAMBDA=0.022,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=1.50E-05,VTO=-0.5,LAMBDA=0.047)
.MODEL NIX NMOS (LEVEL=2,KP=4.00E-05,VTO=0.5,LAMBDA=0.022)
.MODEL DX D(IS=1E-14,RS=5)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=4.84E-11)
*
*
.ENDS AD8617





